`include "mux_dataflow.v"


module mux(in, sel, out);
	input [7:0] in;
	input [2:0]sel;
	output out;
mux
	endmodule 
