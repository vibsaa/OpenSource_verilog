module test();


