module sub32(a,b,sub);
input [31:0]a ,b;
output [31:0] sub;

assign sub=a-b;

endmodule
