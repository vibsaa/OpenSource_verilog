module test();

wire valid;
reg addr;
reg [32:0] wdata;
reg [63:1] rdata;
wire [7:0] write_data;

endmodule
