module mul16(p,q,r);
//how to do this one becuase if both inputs are of 32 widht then result would be so large and require more than 32 bits



endmodule
